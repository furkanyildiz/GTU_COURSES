library verilog;
use verilog.vl_types.all;
entity like_alu_testbench is
end like_alu_testbench;
