module five_bit_and_gate(out,inpA,inpB);

input inpA, inpB;
output out ;
wire out;

endmodule